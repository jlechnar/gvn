../verilog/halve_adder.v