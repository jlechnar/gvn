../verilog/full_adder.v