../verilog/carry_ripple_adder.v